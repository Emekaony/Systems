// this is hello world example
module hello_world();
    // display the message
    initial begin
        $display("Hellow world"); // turns out I don't even need the newline
        $display("Emeka really out here writing verilog huh");
    end
endmodule